`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/05/23 18:22:12
// Design Name: 
// Module Name: PC
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC(
input clk,
input rst,
input PC_W,
input [31:0] data_in,
output reg [31:0] data_out
    );
always @(posedge clk, posedge rst)
begin
if (rst)
    data_out <= 32'b0;
else if (PC_W)
    data_out <= data_in;
else
    data_out <= data_out;
end

endmodule
